// image_parallel_processing_qsys_proc_0_0.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module image_parallel_processing_qsys_proc_0_0 (
		input  wire        clk_clk,                         //               clk.clk
		input  wire        out_bridge_master_waitrequest,   // out_bridge_master.waitrequest
		input  wire [31:0] out_bridge_master_readdata,      //                  .readdata
		input  wire        out_bridge_master_readdatavalid, //                  .readdatavalid
		output wire [0:0]  out_bridge_master_burstcount,    //                  .burstcount
		output wire [31:0] out_bridge_master_writedata,     //                  .writedata
		output wire [26:0] out_bridge_master_address,       //                  .address
		output wire        out_bridge_master_write,         //                  .write
		output wire        out_bridge_master_read,          //                  .read
		output wire [3:0]  out_bridge_master_byteenable,    //                  .byteenable
		output wire        out_bridge_master_debugaccess,   //                  .debugaccess
		input  wire        reset_reset_n                    //             reset.reset_n
	);

	wire  [31:0] proc_0_data_master_readdata;                                 // mm_interconnect_0:proc_0_data_master_readdata -> proc_0:d_readdata
	wire         proc_0_data_master_waitrequest;                              // mm_interconnect_0:proc_0_data_master_waitrequest -> proc_0:d_waitrequest
	wire         proc_0_data_master_debugaccess;                              // proc_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:proc_0_data_master_debugaccess
	wire  [27:0] proc_0_data_master_address;                                  // proc_0:d_address -> mm_interconnect_0:proc_0_data_master_address
	wire   [3:0] proc_0_data_master_byteenable;                               // proc_0:d_byteenable -> mm_interconnect_0:proc_0_data_master_byteenable
	wire         proc_0_data_master_read;                                     // proc_0:d_read -> mm_interconnect_0:proc_0_data_master_read
	wire         proc_0_data_master_readdatavalid;                            // mm_interconnect_0:proc_0_data_master_readdatavalid -> proc_0:d_readdatavalid
	wire         proc_0_data_master_write;                                    // proc_0:d_write -> mm_interconnect_0:proc_0_data_master_write
	wire  [31:0] proc_0_data_master_writedata;                                // proc_0:d_writedata -> mm_interconnect_0:proc_0_data_master_writedata
	wire  [31:0] proc_0_instruction_master_readdata;                          // mm_interconnect_0:proc_0_instruction_master_readdata -> proc_0:i_readdata
	wire         proc_0_instruction_master_waitrequest;                       // mm_interconnect_0:proc_0_instruction_master_waitrequest -> proc_0:i_waitrequest
	wire  [16:0] proc_0_instruction_master_address;                           // proc_0:i_address -> mm_interconnect_0:proc_0_instruction_master_address
	wire         proc_0_instruction_master_read;                              // proc_0:i_read -> mm_interconnect_0:proc_0_instruction_master_read
	wire         proc_0_instruction_master_readdatavalid;                     // mm_interconnect_0:proc_0_instruction_master_readdatavalid -> proc_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_proc_0_debug_mem_slave_readdata;           // proc_0:debug_mem_slave_readdata -> mm_interconnect_0:proc_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_proc_0_debug_mem_slave_waitrequest;        // proc_0:debug_mem_slave_waitrequest -> mm_interconnect_0:proc_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_proc_0_debug_mem_slave_debugaccess;        // mm_interconnect_0:proc_0_debug_mem_slave_debugaccess -> proc_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_proc_0_debug_mem_slave_address;            // mm_interconnect_0:proc_0_debug_mem_slave_address -> proc_0:debug_mem_slave_address
	wire         mm_interconnect_0_proc_0_debug_mem_slave_read;               // mm_interconnect_0:proc_0_debug_mem_slave_read -> proc_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_proc_0_debug_mem_slave_byteenable;         // mm_interconnect_0:proc_0_debug_mem_slave_byteenable -> proc_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_proc_0_debug_mem_slave_write;              // mm_interconnect_0:proc_0_debug_mem_slave_write -> proc_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_proc_0_debug_mem_slave_writedata;          // mm_interconnect_0:proc_0_debug_mem_slave_writedata -> proc_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_out_bridg_0_s0_readdata;                   // out_bridg_0:s0_readdata -> mm_interconnect_0:out_bridg_0_s0_readdata
	wire         mm_interconnect_0_out_bridg_0_s0_waitrequest;                // out_bridg_0:s0_waitrequest -> mm_interconnect_0:out_bridg_0_s0_waitrequest
	wire         mm_interconnect_0_out_bridg_0_s0_debugaccess;                // mm_interconnect_0:out_bridg_0_s0_debugaccess -> out_bridg_0:s0_debugaccess
	wire  [26:0] mm_interconnect_0_out_bridg_0_s0_address;                    // mm_interconnect_0:out_bridg_0_s0_address -> out_bridg_0:s0_address
	wire         mm_interconnect_0_out_bridg_0_s0_read;                       // mm_interconnect_0:out_bridg_0_s0_read -> out_bridg_0:s0_read
	wire   [3:0] mm_interconnect_0_out_bridg_0_s0_byteenable;                 // mm_interconnect_0:out_bridg_0_s0_byteenable -> out_bridg_0:s0_byteenable
	wire         mm_interconnect_0_out_bridg_0_s0_readdatavalid;              // out_bridg_0:s0_readdatavalid -> mm_interconnect_0:out_bridg_0_s0_readdatavalid
	wire         mm_interconnect_0_out_bridg_0_s0_write;                      // mm_interconnect_0:out_bridg_0_s0_write -> out_bridg_0:s0_write
	wire  [31:0] mm_interconnect_0_out_bridg_0_s0_writedata;                  // mm_interconnect_0:out_bridg_0_s0_writedata -> out_bridg_0:s0_writedata
	wire   [0:0] mm_interconnect_0_out_bridg_0_s0_burstcount;                 // mm_interconnect_0:out_bridg_0_s0_burstcount -> out_bridg_0:s0_burstcount
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] proc_0_irq_irq;                                              // irq_mapper:sender_irq -> proc_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:proc_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, out_bridg_0:reset, proc_0:reset_n, rst_translator:in_reset, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [onchip_memory2_0:reset_req, proc_0:reset_req, rst_translator:reset_req_in]

	image_parallel_processing_qsys_proc_0_0_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	image_parallel_processing_qsys_proc_0_0_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (27),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) out_bridg_0 (
		.clk              (clk_clk),                                        //   clk.clk
		.reset            (rst_controller_reset_out_reset),                 // reset.reset
		.s0_waitrequest   (mm_interconnect_0_out_bridg_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_out_bridg_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_out_bridg_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_out_bridg_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_out_bridg_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_out_bridg_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_out_bridg_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_out_bridg_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_out_bridg_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_out_bridg_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (out_bridge_master_waitrequest),                  //    m0.waitrequest
		.m0_readdata      (out_bridge_master_readdata),                     //      .readdata
		.m0_readdatavalid (out_bridge_master_readdatavalid),                //      .readdatavalid
		.m0_burstcount    (out_bridge_master_burstcount),                   //      .burstcount
		.m0_writedata     (out_bridge_master_writedata),                    //      .writedata
		.m0_address       (out_bridge_master_address),                      //      .address
		.m0_write         (out_bridge_master_write),                        //      .write
		.m0_read          (out_bridge_master_read),                         //      .read
		.m0_byteenable    (out_bridge_master_byteenable),                   //      .byteenable
		.m0_debugaccess   (out_bridge_master_debugaccess),                  //      .debugaccess
		.s0_response      (),                                               // (terminated)
		.m0_response      (2'b00)                                           // (terminated)
	);

	image_parallel_processing_qsys_proc_0_0_proc_0 proc_0 (
		.clk                                 (clk_clk),                                              //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (proc_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (proc_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (proc_0_data_master_read),                              //                          .read
		.d_readdata                          (proc_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (proc_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (proc_0_data_master_write),                             //                          .write
		.d_writedata                         (proc_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (proc_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (proc_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (proc_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (proc_0_instruction_master_read),                       //                          .read
		.i_readdata                          (proc_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (proc_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (proc_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (proc_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_proc_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_proc_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_proc_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_proc_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_proc_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_proc_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_proc_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_proc_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	image_parallel_processing_qsys_proc_0_0_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	image_parallel_processing_qsys_proc_0_0_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                             (clk_clk),                                                     //                          clk_0_clk.clk
		.proc_0_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                              // proc_0_reset_reset_bridge_in_reset.reset
		.proc_0_data_master_address                (proc_0_data_master_address),                                  //                 proc_0_data_master.address
		.proc_0_data_master_waitrequest            (proc_0_data_master_waitrequest),                              //                                   .waitrequest
		.proc_0_data_master_byteenable             (proc_0_data_master_byteenable),                               //                                   .byteenable
		.proc_0_data_master_read                   (proc_0_data_master_read),                                     //                                   .read
		.proc_0_data_master_readdata               (proc_0_data_master_readdata),                                 //                                   .readdata
		.proc_0_data_master_readdatavalid          (proc_0_data_master_readdatavalid),                            //                                   .readdatavalid
		.proc_0_data_master_write                  (proc_0_data_master_write),                                    //                                   .write
		.proc_0_data_master_writedata              (proc_0_data_master_writedata),                                //                                   .writedata
		.proc_0_data_master_debugaccess            (proc_0_data_master_debugaccess),                              //                                   .debugaccess
		.proc_0_instruction_master_address         (proc_0_instruction_master_address),                           //          proc_0_instruction_master.address
		.proc_0_instruction_master_waitrequest     (proc_0_instruction_master_waitrequest),                       //                                   .waitrequest
		.proc_0_instruction_master_read            (proc_0_instruction_master_read),                              //                                   .read
		.proc_0_instruction_master_readdata        (proc_0_instruction_master_readdata),                          //                                   .readdata
		.proc_0_instruction_master_readdatavalid   (proc_0_instruction_master_readdatavalid),                     //                                   .readdatavalid
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //      jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                   .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                   .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                   .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                   .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                   .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                   .chipselect
		.onchip_memory2_0_s1_address               (mm_interconnect_0_onchip_memory2_0_s1_address),               //                onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                 (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                   .write
		.onchip_memory2_0_s1_readdata              (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                   .readdata
		.onchip_memory2_0_s1_writedata             (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                   .writedata
		.onchip_memory2_0_s1_byteenable            (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                   .byteenable
		.onchip_memory2_0_s1_chipselect            (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                   .chipselect
		.onchip_memory2_0_s1_clken                 (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                   .clken
		.out_bridg_0_s0_address                    (mm_interconnect_0_out_bridg_0_s0_address),                    //                     out_bridg_0_s0.address
		.out_bridg_0_s0_write                      (mm_interconnect_0_out_bridg_0_s0_write),                      //                                   .write
		.out_bridg_0_s0_read                       (mm_interconnect_0_out_bridg_0_s0_read),                       //                                   .read
		.out_bridg_0_s0_readdata                   (mm_interconnect_0_out_bridg_0_s0_readdata),                   //                                   .readdata
		.out_bridg_0_s0_writedata                  (mm_interconnect_0_out_bridg_0_s0_writedata),                  //                                   .writedata
		.out_bridg_0_s0_burstcount                 (mm_interconnect_0_out_bridg_0_s0_burstcount),                 //                                   .burstcount
		.out_bridg_0_s0_byteenable                 (mm_interconnect_0_out_bridg_0_s0_byteenable),                 //                                   .byteenable
		.out_bridg_0_s0_readdatavalid              (mm_interconnect_0_out_bridg_0_s0_readdatavalid),              //                                   .readdatavalid
		.out_bridg_0_s0_waitrequest                (mm_interconnect_0_out_bridg_0_s0_waitrequest),                //                                   .waitrequest
		.out_bridg_0_s0_debugaccess                (mm_interconnect_0_out_bridg_0_s0_debugaccess),                //                                   .debugaccess
		.proc_0_debug_mem_slave_address            (mm_interconnect_0_proc_0_debug_mem_slave_address),            //             proc_0_debug_mem_slave.address
		.proc_0_debug_mem_slave_write              (mm_interconnect_0_proc_0_debug_mem_slave_write),              //                                   .write
		.proc_0_debug_mem_slave_read               (mm_interconnect_0_proc_0_debug_mem_slave_read),               //                                   .read
		.proc_0_debug_mem_slave_readdata           (mm_interconnect_0_proc_0_debug_mem_slave_readdata),           //                                   .readdata
		.proc_0_debug_mem_slave_writedata          (mm_interconnect_0_proc_0_debug_mem_slave_writedata),          //                                   .writedata
		.proc_0_debug_mem_slave_byteenable         (mm_interconnect_0_proc_0_debug_mem_slave_byteenable),         //                                   .byteenable
		.proc_0_debug_mem_slave_waitrequest        (mm_interconnect_0_proc_0_debug_mem_slave_waitrequest),        //                                   .waitrequest
		.proc_0_debug_mem_slave_debugaccess        (mm_interconnect_0_proc_0_debug_mem_slave_debugaccess),        //                                   .debugaccess
		.timer_0_s1_address                        (mm_interconnect_0_timer_0_s1_address),                        //                         timer_0_s1.address
		.timer_0_s1_write                          (mm_interconnect_0_timer_0_s1_write),                          //                                   .write
		.timer_0_s1_readdata                       (mm_interconnect_0_timer_0_s1_readdata),                       //                                   .readdata
		.timer_0_s1_writedata                      (mm_interconnect_0_timer_0_s1_writedata),                      //                                   .writedata
		.timer_0_s1_chipselect                     (mm_interconnect_0_timer_0_s1_chipselect)                      //                                   .chipselect
	);

	image_parallel_processing_qsys_proc_0_0_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (proc_0_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
